`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Hextio Inc.
// Engineer: Kamil KAYA
// 
// Create Date:    14:37:28 10/22/2018 
// Design Name: 	 UART HARDWARE DESIGN
// Module Name:    UART Receive Module
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
//--------------------------------------------------------------------------------
module UART_RX(input SYSCLK,
				input [7:0] DATA,
				input SEND,
				output reg BUSY_FLAG,
				output reg COMPLATE_FLAG,
				output reg ERROR_FLAG);



endmodule
