`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 	
// Engineer: 	Kamil KAYA
// 
// Create Date: 02/13/2021 07:33:04 PM
// Design Name: 
// Module Name: And Gate
// Project Name: 	Tutorial
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module andgate(input a, input b, output q);

assign q=a & b;

endmodule
